Library IEEE;
Use IEEE.std_logic_1164.all;
Use IEEE.std_logic_unsigned.all;
----------------------------------------
entity basic_structure is
	port(
	
	);
end basic_structure;
-----------------------------------------
architecture test1 of basic_structure is
	
begin
	process()
	
	begin
	
	end process;
end test1;











