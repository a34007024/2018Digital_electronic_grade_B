Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logoc_unsigned.all;

entity nox1_180810 is
	port();
	
end entity;

architecture main of nox1_180810 is

begin

end architecture;