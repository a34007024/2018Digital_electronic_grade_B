Library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
----------------------------------
Entity Nox1_practice is

End Nox1_practice;